module cnt_cam
#(
  parameter CNT_SIZE    = 13, /*tbd*/ 
  parameter NUM_ENTRY   = 50,
  parameter ENTRY_WIDTH = 6, // [log2(NUM_ENTRY)]
  parameter TOP_K       = 5
)
(
  input                    clk,
  input                    reset,
  input                    incremental_en,
  input                    sort_en,
  input                    mig_en,
  input  [ENTRY_WIDTH-1:0] incremental_rank,
  input  [ENTRY_WIDTH-1:0] hit_compare_rank,
  input  [ENTRY_WIDTH-1:0] sort_hit_rank,
  input  [ENTRY_WIDTH-1:0] minptr,
  output [ENTRY_WIDTH-1:0] new_minptr,
  output [ENTRY_WIDTH-1:0] new_rank,
  output [CNT_SIZE-1:0]    top_1,
  output [CNT_SIZE-1:0]    top_2,
  output [CNT_SIZE-1:0]    top_3,
  output [CNT_SIZE-1:0]    top_4,
  output [CNT_SIZE-1:0]    top_5,
  input  [2:0]             num_mig
);

  wire                   we_array             [0:NUM_ENTRY-1];
  wire [CNT_SIZE-1:0]    data_array_in        [0:NUM_ENTRY-1];

  reg  [CNT_SIZE-1:0]    sort_data_array_in   [0:NUM_ENTRY-1];
  reg  [CNT_SIZE-1:0]    mig_data_array_in    [0:NUM_ENTRY-1];

  wire [CNT_SIZE-1:0]    data_array_out       [0:NUM_ENTRY-1];
  wire [CNT_SIZE-1:0]    hit_refer;
  wire [CNT_SIZE-1:0]    miss_refer;
  reg  [NUM_ENTRY-1:0]   hit_compare_result;
  reg  [NUM_ENTRY-1:0]   miss_compare_result;

  reg  [ENTRY_WIDTH:0]   hit_zeros;
  reg  [ENTRY_WIDTH:0]   miss_zeros;

  reg  [ENTRY_WIDTH-1:0] new_minptr_r;

  wire                   top_k_cache_table_we;
  wire [CNT_SIZE-1:0]    top_k_data_array_in  [0:TOP_K-1];
  wire [CNT_SIZE-1:0]    top_k_data_array_out [0:TOP_K-1];


  genvar i, j, k;
  integer h;

  generate for (i = 0; i < NUM_ENTRY; i = i+1) begin: ffarray_inst
      assign we_array[i]      = reset ? 1 : ((incremental_en & (incremental_rank == i)) || sort_en || mig_en);
      assign data_array_in[i] = reset ? 0 :
                                        incremental_en ? (data_array_out[i] + 1) : 
                                                         sort_en ? sort_data_array_in[i] :
                                                                   mig_en ? mig_data_array_in[i] :
                                                                            0;

      FF_array
      #(
        .WORD_SIZE ( CNT_SIZE )
      )
        FF_array_
      (
        .clk       ( clk               ),
        .data_in   ( data_array_in[i]  ),
        .write_en  ( we_array[i]       ),
        .search_en ( 1'b0              ),
        .data_out  ( data_array_out[i] ),
        .match     (                   )
      );
  end
  endgenerate


  generate for (j = 0; j < NUM_ENTRY; j = j + 1) begin
      always_comb begin   
        if (sort_en) begin
          if(j == new_rank) begin
            sort_data_array_in[j] = data_array_out[sort_hit_rank] + 1;
          end
          else if ((j <= sort_hit_rank) && (j > new_rank)) begin
            sort_data_array_in[j] = data_array_out[j-1];
          end 
          else begin
            sort_data_array_in[j] = data_array_out[j];
          end
        end
        else begin
          sort_data_array_in[j] = 0;
        end
      end

      always_comb begin   
        if (mig_en & (j <= NUM_ENTRY - 1 - num_mig)) begin
          mig_data_array_in[j] = data_array_out[j+num_mig] - data_array_out[minptr];
        end
        else begin
          mig_data_array_in[j] = 0;
        end
      end
  end
  endgenerate


  assign hit_refer = data_array_out[hit_compare_rank];
  assign miss_refer = data_array_out[minptr]+1;

  // when hit or miss_compare_en, compare CAM's count value with (hit rank's count+1) or (minptr_count + 1) 
  generate for (k = 0; k < NUM_ENTRY; k = k+1) begin
    always_ff @(posedge clk or posedge reset) begin
      if (reset) begin
        hit_compare_result[k] <= 0;
        miss_compare_result[k] <= 0;
      end
      else begin
        hit_compare_result[k] <= (hit_refer >= data_array_out[k]);
        miss_compare_result[k] <= (miss_refer >= data_array_out[k]);
      end
    end
  end
  endgenerate

  /*
  always_comb begin
    case(hit_compare_result)
      100'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd99;
      100'b1100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd98;
      100'b1110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd97;
      100'b1111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd96;
      100'b1111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd95;
      100'b1111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd94;
      100'b1111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd93;
      100'b1111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd92;
      100'b1111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd91;
      100'b1111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd90;
      100'b1111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd89;
      100'b1111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd88;
      100'b1111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd87;
      100'b1111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd86;
      100'b1111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd85;
      100'b1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd84;
      100'b1111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd83;
      100'b1111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd82;
      100'b1111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd81;
      100'b1111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd80;
      100'b1111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd79;
      100'b1111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd78;
      100'b1111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd77;
      100'b1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd76;
      100'b1111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd75;
      100'b1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd74;
      100'b1111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd73;
      100'b1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd72;
      100'b1111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd71;
      100'b1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd70;
      100'b1111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd69;
      100'b1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd68;
      100'b1111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd67;
      100'b1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd66;
      100'b1111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd65;
      100'b1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd64;
      100'b1111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd63;
      100'b1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd62;
      100'b1111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd61;
      100'b1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd60;
      100'b1111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd59;
      100'b1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd58;
      100'b1111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd57;
      100'b1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd56;
      100'b1111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd55;
      100'b1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000: hit_zeros = 7'd54;
      100'b1111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000: hit_zeros = 7'd53;
      100'b1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000: hit_zeros = 7'd52;
      100'b1111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000: hit_zeros = 7'd51;
      100'b1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000: hit_zeros = 7'd50;
      100'b1111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000: hit_zeros = 7'd49;
      100'b1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000: hit_zeros = 7'd48;
      100'b1111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000: hit_zeros = 7'd47;
      100'b1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000: hit_zeros = 7'd46;
      100'b1111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000: hit_zeros = 7'd45;
      100'b1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000: hit_zeros = 7'd44;
      100'b1111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000: hit_zeros = 7'd43;
      100'b1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000: hit_zeros = 7'd42;
      100'b1111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000: hit_zeros = 7'd41;
      100'b1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000: hit_zeros = 7'd40;
      100'b1111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000: hit_zeros = 7'd39;
      100'b1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000: hit_zeros = 7'd38;
      100'b1111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000: hit_zeros = 7'd37;
      100'b1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000: hit_zeros = 7'd36;
      100'b1111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000: hit_zeros = 7'd35;
      100'b1111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000: hit_zeros = 7'd34;
      100'b1111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000: hit_zeros = 7'd33;
      100'b1111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000: hit_zeros = 7'd32;
      100'b1111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000: hit_zeros = 7'd31;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000: hit_zeros = 7'd30;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000: hit_zeros = 7'd29;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000: hit_zeros = 7'd28;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000: hit_zeros = 7'd27;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000: hit_zeros = 7'd26;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000: hit_zeros = 7'd25;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000: hit_zeros = 7'd24;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000: hit_zeros = 7'd23;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000: hit_zeros = 7'd22;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000: hit_zeros = 7'd21;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000: hit_zeros = 7'd20;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000: hit_zeros = 7'd19;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000: hit_zeros = 7'd18;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000: hit_zeros = 7'd17;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000: hit_zeros = 7'd16;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000: hit_zeros = 7'd15;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000: hit_zeros = 7'd14;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000: hit_zeros = 7'd13;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000: hit_zeros = 7'd12;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000: hit_zeros = 7'd11;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000: hit_zeros = 7'd10;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000: hit_zeros = 7'd9;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000: hit_zeros = 7'd8;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000: hit_zeros = 7'd7;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000: hit_zeros = 7'd6;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000: hit_zeros = 7'd5;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000: hit_zeros = 7'd4;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000: hit_zeros = 7'd3;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100: hit_zeros = 7'd2;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110: hit_zeros = 7'd1;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: hit_zeros = 7'd0;
      default: hit_zeros = 7'd0;
    endcase
  end
  always_comb begin
    case(miss_compare_result)
      100'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd99;
      100'b1100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd98;
      100'b1110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd97;
      100'b1111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd96;
      100'b1111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd95;
      100'b1111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd94;
      100'b1111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd93;
      100'b1111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd92;
      100'b1111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd91;
      100'b1111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd90;
      100'b1111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd89;
      100'b1111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd88;
      100'b1111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd87;
      100'b1111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd86;
      100'b1111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd85;
      100'b1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd84;
      100'b1111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd83;
      100'b1111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd82;
      100'b1111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd81;
      100'b1111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd80;
      100'b1111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd79;
      100'b1111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd78;
      100'b1111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd77;
      100'b1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd76;
      100'b1111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd75;
      100'b1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd74;
      100'b1111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd73;
      100'b1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd72;
      100'b1111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd71;
      100'b1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd70;
      100'b1111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd69;
      100'b1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd68;
      100'b1111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd67;
      100'b1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd66;
      100'b1111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd65;
      100'b1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd64;
      100'b1111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd63;
      100'b1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd62;
      100'b1111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd61;
      100'b1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd60;
      100'b1111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd59;
      100'b1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd58;
      100'b1111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd57;
      100'b1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd56;
      100'b1111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd55;
      100'b1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000: miss_zeros = 7'd54;
      100'b1111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000: miss_zeros = 7'd53;
      100'b1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000: miss_zeros = 7'd52;
      100'b1111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000: miss_zeros = 7'd51;
      100'b1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000: miss_zeros = 7'd50;
      100'b1111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000: miss_zeros = 7'd49;
      100'b1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000: miss_zeros = 7'd48;
      100'b1111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000: miss_zeros = 7'd47;
      100'b1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000: miss_zeros = 7'd46;
      100'b1111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000: miss_zeros = 7'd45;
      100'b1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000: miss_zeros = 7'd44;
      100'b1111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000: miss_zeros = 7'd43;
      100'b1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000: miss_zeros = 7'd42;
      100'b1111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000: miss_zeros = 7'd41;
      100'b1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000: miss_zeros = 7'd40;
      100'b1111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000: miss_zeros = 7'd39;
      100'b1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000: miss_zeros = 7'd38;
      100'b1111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000: miss_zeros = 7'd37;
      100'b1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000: miss_zeros = 7'd36;
      100'b1111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000: miss_zeros = 7'd35;
      100'b1111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000: miss_zeros = 7'd34;
      100'b1111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000: miss_zeros = 7'd33;
      100'b1111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000: miss_zeros = 7'd32;
      100'b1111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000: miss_zeros = 7'd31;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000: miss_zeros = 7'd30;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000: miss_zeros = 7'd29;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000: miss_zeros = 7'd28;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000: miss_zeros = 7'd27;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000: miss_zeros = 7'd26;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000: miss_zeros = 7'd25;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000: miss_zeros = 7'd24;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000: miss_zeros = 7'd23;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000: miss_zeros = 7'd22;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000: miss_zeros = 7'd21;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000: miss_zeros = 7'd20;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000: miss_zeros = 7'd19;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000: miss_zeros = 7'd18;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000: miss_zeros = 7'd17;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000: miss_zeros = 7'd16;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000: miss_zeros = 7'd15;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000: miss_zeros = 7'd14;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000: miss_zeros = 7'd13;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000: miss_zeros = 7'd12;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000: miss_zeros = 7'd11;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000: miss_zeros = 7'd10;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000: miss_zeros = 7'd9;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000: miss_zeros = 7'd8;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000: miss_zeros = 7'd7;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000: miss_zeros = 7'd6;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000: miss_zeros = 7'd5;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000: miss_zeros = 7'd4;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000: miss_zeros = 7'd3;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100: miss_zeros = 7'd2;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110: miss_zeros = 7'd1;
      100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: miss_zeros = 7'd0;
      default: miss_zeros = 7'd0;
    endcase
  end
  */


  always_comb begin
    case(hit_compare_result)
      50'b10000000000000000000000000000000000000000000000000: hit_zeros = 6'd49;
      50'b11000000000000000000000000000000000000000000000000: hit_zeros = 6'd48;
      50'b11100000000000000000000000000000000000000000000000: hit_zeros = 6'd47;
      50'b11110000000000000000000000000000000000000000000000: hit_zeros = 6'd46;
      50'b11111000000000000000000000000000000000000000000000: hit_zeros = 6'd45;
      50'b11111100000000000000000000000000000000000000000000: hit_zeros = 6'd44;
      50'b11111110000000000000000000000000000000000000000000: hit_zeros = 6'd43;
      50'b11111111000000000000000000000000000000000000000000: hit_zeros = 6'd42;
      50'b11111111100000000000000000000000000000000000000000: hit_zeros = 6'd41;
      50'b11111111110000000000000000000000000000000000000000: hit_zeros = 6'd40;
      50'b11111111111000000000000000000000000000000000000000: hit_zeros = 6'd39;
      50'b11111111111100000000000000000000000000000000000000: hit_zeros = 6'd38;
      50'b11111111111110000000000000000000000000000000000000: hit_zeros = 6'd37;
      50'b11111111111111000000000000000000000000000000000000: hit_zeros = 6'd36;
      50'b11111111111111100000000000000000000000000000000000: hit_zeros = 6'd35;
      50'b11111111111111110000000000000000000000000000000000: hit_zeros = 6'd34;
      50'b11111111111111111000000000000000000000000000000000: hit_zeros = 6'd33;
      50'b11111111111111111100000000000000000000000000000000: hit_zeros = 6'd32;
      50'b11111111111111111110000000000000000000000000000000: hit_zeros = 6'd31;
      50'b11111111111111111111000000000000000000000000000000: hit_zeros = 6'd30;
      50'b11111111111111111111100000000000000000000000000000: hit_zeros = 6'd29;
      50'b11111111111111111111110000000000000000000000000000: hit_zeros = 6'd28;
      50'b11111111111111111111111000000000000000000000000000: hit_zeros = 6'd27;
      50'b11111111111111111111111100000000000000000000000000: hit_zeros = 6'd26;
      50'b11111111111111111111111110000000000000000000000000: hit_zeros = 6'd25;
      50'b11111111111111111111111111000000000000000000000000: hit_zeros = 6'd24;
      50'b11111111111111111111111111100000000000000000000000: hit_zeros = 6'd23;
      50'b11111111111111111111111111110000000000000000000000: hit_zeros = 6'd22;
      50'b11111111111111111111111111111000000000000000000000: hit_zeros = 6'd21;
      50'b11111111111111111111111111111100000000000000000000: hit_zeros = 6'd20;
      50'b11111111111111111111111111111110000000000000000000: hit_zeros = 6'd19;
      50'b11111111111111111111111111111111000000000000000000: hit_zeros = 6'd18;
      50'b11111111111111111111111111111111100000000000000000: hit_zeros = 6'd17;
      50'b11111111111111111111111111111111110000000000000000: hit_zeros = 6'd16;
      50'b11111111111111111111111111111111111000000000000000: hit_zeros = 6'd15;
      50'b11111111111111111111111111111111111100000000000000: hit_zeros = 6'd14;
      50'b11111111111111111111111111111111111110000000000000: hit_zeros = 6'd13;
      50'b11111111111111111111111111111111111111000000000000: hit_zeros = 6'd12;
      50'b11111111111111111111111111111111111111100000000000: hit_zeros = 6'd11;
      50'b11111111111111111111111111111111111111110000000000: hit_zeros = 6'd10;
      50'b11111111111111111111111111111111111111111000000000: hit_zeros = 6'd9;
      50'b11111111111111111111111111111111111111111100000000: hit_zeros = 6'd8;
      50'b11111111111111111111111111111111111111111110000000: hit_zeros = 6'd7;
      50'b11111111111111111111111111111111111111111111000000: hit_zeros = 6'd6;
      50'b11111111111111111111111111111111111111111111100000: hit_zeros = 6'd5;
      50'b11111111111111111111111111111111111111111111110000: hit_zeros = 6'd4;
      50'b11111111111111111111111111111111111111111111111000: hit_zeros = 6'd3;
      50'b11111111111111111111111111111111111111111111111100: hit_zeros = 6'd2;
      50'b11111111111111111111111111111111111111111111111110: hit_zeros = 6'd1;
      50'b11111111111111111111111111111111111111111111111111: hit_zeros = 6'd0;
      default: hit_zeros = 7'd0;
    endcase
  end
  always_comb begin
    case(miss_compare_result)
      50'b10000000000000000000000000000000000000000000000000: miss_zeros = 6'd49;
      50'b11000000000000000000000000000000000000000000000000: miss_zeros = 6'd48;
      50'b11100000000000000000000000000000000000000000000000: miss_zeros = 6'd47;
      50'b11110000000000000000000000000000000000000000000000: miss_zeros = 6'd46;
      50'b11111000000000000000000000000000000000000000000000: miss_zeros = 6'd45;
      50'b11111100000000000000000000000000000000000000000000: miss_zeros = 6'd44;
      50'b11111110000000000000000000000000000000000000000000: miss_zeros = 6'd43;
      50'b11111111000000000000000000000000000000000000000000: miss_zeros = 6'd42;
      50'b11111111100000000000000000000000000000000000000000: miss_zeros = 6'd41;
      50'b11111111110000000000000000000000000000000000000000: miss_zeros = 6'd40;
      50'b11111111111000000000000000000000000000000000000000: miss_zeros = 6'd39;
      50'b11111111111100000000000000000000000000000000000000: miss_zeros = 6'd38;
      50'b11111111111110000000000000000000000000000000000000: miss_zeros = 6'd37;
      50'b11111111111111000000000000000000000000000000000000: miss_zeros = 6'd36;
      50'b11111111111111100000000000000000000000000000000000: miss_zeros = 6'd35;
      50'b11111111111111110000000000000000000000000000000000: miss_zeros = 6'd34;
      50'b11111111111111111000000000000000000000000000000000: miss_zeros = 6'd33;
      50'b11111111111111111100000000000000000000000000000000: miss_zeros = 6'd32;
      50'b11111111111111111110000000000000000000000000000000: miss_zeros = 6'd31;
      50'b11111111111111111111000000000000000000000000000000: miss_zeros = 6'd30;
      50'b11111111111111111111100000000000000000000000000000: miss_zeros = 6'd29;
      50'b11111111111111111111110000000000000000000000000000: miss_zeros = 6'd28;
      50'b11111111111111111111111000000000000000000000000000: miss_zeros = 6'd27;
      50'b11111111111111111111111100000000000000000000000000: miss_zeros = 6'd26;
      50'b11111111111111111111111110000000000000000000000000: miss_zeros = 6'd25;
      50'b11111111111111111111111111000000000000000000000000: miss_zeros = 6'd24;
      50'b11111111111111111111111111100000000000000000000000: miss_zeros = 6'd23;
      50'b11111111111111111111111111110000000000000000000000: miss_zeros = 6'd22;
      50'b11111111111111111111111111111000000000000000000000: miss_zeros = 6'd21;
      50'b11111111111111111111111111111100000000000000000000: miss_zeros = 6'd20;
      50'b11111111111111111111111111111110000000000000000000: miss_zeros = 6'd19;
      50'b11111111111111111111111111111111000000000000000000: miss_zeros = 6'd18;
      50'b11111111111111111111111111111111100000000000000000: miss_zeros = 6'd17;
      50'b11111111111111111111111111111111110000000000000000: miss_zeros = 6'd16;
      50'b11111111111111111111111111111111111000000000000000: miss_zeros = 6'd15;
      50'b11111111111111111111111111111111111100000000000000: miss_zeros = 6'd14;
      50'b11111111111111111111111111111111111110000000000000: miss_zeros = 6'd13;
      50'b11111111111111111111111111111111111111000000000000: miss_zeros = 6'd12;
      50'b11111111111111111111111111111111111111100000000000: miss_zeros = 6'd11;
      50'b11111111111111111111111111111111111111110000000000: miss_zeros = 6'd10;
      50'b11111111111111111111111111111111111111111000000000: miss_zeros = 6'd9;
      50'b11111111111111111111111111111111111111111100000000: miss_zeros = 6'd8;
      50'b11111111111111111111111111111111111111111110000000: miss_zeros = 6'd7;
      50'b11111111111111111111111111111111111111111111000000: miss_zeros = 6'd6;
      50'b11111111111111111111111111111111111111111111100000: miss_zeros = 6'd5;
      50'b11111111111111111111111111111111111111111111110000: miss_zeros = 6'd4;
      50'b11111111111111111111111111111111111111111111111000: miss_zeros = 6'd3;
      50'b11111111111111111111111111111111111111111111111100: miss_zeros = 6'd2;
      50'b11111111111111111111111111111111111111111111111110: miss_zeros = 6'd1;
      50'b11111111111111111111111111111111111111111111111111: miss_zeros = 6'd0;
      default: miss_zeros = 6'd0;
    endcase
  end

  /*
  // accumulate compare result's number of 1s
  always_comb begin
    hit_zeros = NUM_ENTRY;
    miss_zeros = NUM_ENTRY;
    for(h = 0; h < NUM_ENTRY; h = h + 1) begin
      hit_zeros -= hit_compare_result[h];
      miss_zeros -= miss_compare_result[h];
    end  
  end
  */


  assign new_rank = hit_zeros;

  always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
      new_minptr_r <= {ENTRY_WIDTH{1'b0}};
    end
    else begin
      if (minptr == (NUM_ENTRY - 1)) begin
        new_minptr_r <= miss_zeros;
      end
      else begin
        new_minptr_r <= new_minptr_r;
      end
    end
  end

  assign new_minptr = new_minptr_r;



  /*
  assign top_k_cache_table_we = reset ? 1 : mig_en;

  generate for (k = 0; k < TOP_K; k = k+1) begin: top_k_cache_table_inst

      assign top_k_data_array_in[k] = reset ? 0 : data_array_out[k];

      FF_array #(.WORD_SIZE(CNT_SIZE)) top_k_cache_table(.clk (clk), .data_in(top_k_data_array_in[k]),
        .write_en(top_k_cache_table_we), .search_en(1'b0), .data_out(top_k_data_array_out[k]), .match());
      end
  endgenerate

  assign top_1 = top_k_data_array_out[0];
  assign top_2 = (TOP_K > 1) ? top_k_data_array_out[1] : {CNT_SIZE{1'b0}};
  assign top_3 = (TOP_K > 2) ? top_k_data_array_out[2] : {CNT_SIZE{1'b0}};
  assign top_4 = (TOP_K > 3) ? top_k_data_array_out[3] : {CNT_SIZE{1'b0}};
  assign top_5 = (TOP_K > 4) ? top_k_data_array_out[4] : {CNT_SIZE{1'b0}};
  */

  assign top_1 = data_array_out[0];
  assign top_2 = (TOP_K > 1) ? data_array_out[1] : {CNT_SIZE{1'b0}};
  assign top_3 = (TOP_K > 2) ? data_array_out[2] : {CNT_SIZE{1'b0}};
  assign top_4 = (TOP_K > 3) ? data_array_out[3] : {CNT_SIZE{1'b0}};
  assign top_5 = (TOP_K > 4) ? data_array_out[4] : {CNT_SIZE{1'b0}};

endmodule
